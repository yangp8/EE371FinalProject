module deadPrint ();
	if(dead) 
endmodule
